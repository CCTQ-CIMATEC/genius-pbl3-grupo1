

`ifndef RISCV_DEFINES
`define RISCV_DEFINES

  `define RISCV_WIDTH 4 
  `define NO_OF_TRANSACTIONS 10

`endif
